library ieee;
use ieee.std_logic_1164.all;
use work.Gates.all;

entity ZNVLG  is
  port (X, Y: in std_logic_vector(3 downto 0); Z,N,V,L,G: out std_logic);
end entity ZNVLG;

architecture Struct of ZNVLG is
--write your code here
end Struct;
